`timescale 1ns / 1ps

//`default_nettype none
module BCD_7_Segment(  // Default net type is a wire
    input wire [3:0] data_in,
    output reg [6:0] seg
);

    always @(*)  // Procedural assignments within
    begin
        case(data_in)  // Active low BCD representation
            0: seg = 7'b1000000;
            1: seg = 7'b1111001;
            2: seg = 7'b0100100;
            3: seg = 7'b0110000;
            4: seg = 7'b0011001;
            5: seg = 7'b0010010;
            6: seg = 7'b0000010;
            7: seg = 7'b1111000;
            8: seg = 7'b0000000;
            9: seg = 7'b0010000;
        endcase
    end
endmodule
